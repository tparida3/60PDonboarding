* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  pfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l = l w = w ad = ad as = as pd = pd ps = ps nrd = nrd nrs = nrs sa = sa sb = sb sd = sd nf = nf
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.32+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.041573+sky130_fd_pr__pfet_01v8_lvt__k2_diff_0'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0'
+ ua = '-2.8863e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_0'
+ ub = '2.9625e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_0'
+ uc = 6.4586e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00265+sky130_fd_pr__pfet_01v8_lvt__u0_diff_0'
+ a0 = '1.3255+sky130_fd_pr__pfet_01v8_lvt__a0_diff_0'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_0'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.25696+sky130_fd_pr__pfet_01v8_lvt__ags_diff_0'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_0'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_0'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_0+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.017768
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.046757
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.61727+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0'
+ kt2 = -0.035779
+ at = 164410.0
+ ute = -0.15885
+ ua1 = 6.4145e-10
+ ub1 = -1.094e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.38+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.041573+sky130_fd_pr__pfet_01v8_lvt__k2_diff_1'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1'
+ ua = '-2.8863e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_1'
+ ub = '2.9625e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_1'
+ uc = 6.4586e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00265+sky130_fd_pr__pfet_01v8_lvt__u0_diff_1'
+ a0 = '1.3662+sky130_fd_pr__pfet_01v8_lvt__a0_diff_1'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_1'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.25696+sky130_fd_pr__pfet_01v8_lvt__ags_diff_1'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_1'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_1'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_1+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0091588
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.024056
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1'
+ kt2 = -0.055045
+ at = 240100.0
+ ute = -0.15426
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.38+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.041573+sky130_fd_pr__pfet_01v8_lvt__k2_diff_2'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2'
+ ua = '-2.9363e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_2'
+ ub = '3.023e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_2'
+ uc = 6.4586e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00264+sky130_fd_pr__pfet_01v8_lvt__u0_diff_2'
+ a0 = '1.4534+sky130_fd_pr__pfet_01v8_lvt__a0_diff_2'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_2'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.25696+sky130_fd_pr__pfet_01v8_lvt__ags_diff_2'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_2'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_2'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_2+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0045794
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.022652
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2'
+ kt2 = -0.055045
+ at = 272010.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -7.1909e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.38+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.037416+sky130_fd_pr__pfet_01v8_lvt__k2_diff_3'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3'
+ ua = '-2.8863e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_3'
+ ub = '2.94e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_3'
+ uc = 6.4586e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00254+sky130_fd_pr__pfet_01v8_lvt__u0_diff_3'
+ a0 = '1.3813+sky130_fd_pr__pfet_01v8_lvt__a0_diff_3'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_3'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15932+sky130_fd_pr__pfet_01v8_lvt__ags_diff_3'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_3'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_3'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_3+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0013922
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.012907
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3'
+ kt2 = -0.055045
+ at = 274260.0
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.285+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.016213+sky130_fd_pr__pfet_01v8_lvt__k2_diff_4'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '86632+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4'
+ ua = '-2.9663e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_4'
+ ub = '3.2651e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_4'
+ uc = 5.6836e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.002915+sky130_fd_pr__pfet_01v8_lvt__u0_diff_4'
+ a0 = '1.1627+sky130_fd_pr__pfet_01v8_lvt__a0_diff_4'
+ keta = '-0.011825+sky130_fd_pr__pfet_01v8_lvt__keta_diff_4'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.25696+sky130_fd_pr__pfet_01v8_lvt__ags_diff_4'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_4'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_4'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_4+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.092154
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.051939
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62756+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4'
+ kt2 = -0.085339
+ at = 23556.0
+ ute = -0.21235
+ ua1 = 7.2317e-10
+ ub1 = -2.3247e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.336+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.032427+sky130_fd_pr__pfet_01v8_lvt__k2_diff_5'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5'
+ ua = '-2.9263e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_5'
+ ub = '3.0425e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_5'
+ uc = 5.6836e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00265+sky130_fd_pr__pfet_01v8_lvt__u0_diff_5'
+ a0 = '1.1627+sky130_fd_pr__pfet_01v8_lvt__a0_diff_5'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_5'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.25696+sky130_fd_pr__pfet_01v8_lvt__ags_diff_5'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_5'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_5'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_5+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.049545
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.061832
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.63828+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5'
+ kt2 = -0.050974
+ at = 60707.0
+ ute = -0.23454
+ ua1 = 8.9635e-10
+ ub1 = -6.3517e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos
* DC IV MOS Parameters
+ lmin = 1.495e-06 lmax = 1.505e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.375+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_6'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6'
+ ua = '-2.8887e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_6'
+ ub = '2.8956e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_6'
+ uc = 5.1181e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0028+sky130_fd_pr__pfet_01v8_lvt__u0_diff_6'
+ a0 = '1.4539+sky130_fd_pr__pfet_01v8_lvt__a0_diff_6'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_6'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.20801+sky130_fd_pr__pfet_01v8_lvt__ags_diff_6'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_6'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_6'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_6+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0080176
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.035435
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6'
+ kt2 = -0.055045
+ at = 218490.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.39+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_7'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7'
+ ua = '-2.782e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_7'
+ ub = '2.9317e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_7'
+ uc = '8.3852e-011+sky130_fd_pr__pfet_01v8_lvt__uc_diff_7'
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0033729+sky130_fd_pr__pfet_01v8_lvt__u0_diff_7'
+ a0 = '1.255+sky130_fd_pr__pfet_01v8_lvt__a0_diff_7'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_7'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.3059+sky130_fd_pr__pfet_01v8_lvt__ags_diff_7'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_7'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_7'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_7+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '3.9645+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.012207
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.055778
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7'
+ kt2 = -0.035779
+ at = 186080.0
+ ute = -0.3758
+ ua1 = 6.4145e-10
+ ub1 = -1.094e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.395e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.395+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_8'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8'
+ ua = '-2.8887e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_8'
+ ub = '2.8956e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_8'
+ uc = 5.1181e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0028+sky130_fd_pr__pfet_01v8_lvt__u0_diff_8'
+ a0 = '1.5171+sky130_fd_pr__pfet_01v8_lvt__a0_diff_8'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_8'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.20801+sky130_fd_pr__pfet_01v8_lvt__ags_diff_8'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_8'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_8'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_8+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0064658
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.04
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8'
+ kt2 = -0.055045
+ at = 240100.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 1.765e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.395+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_9'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9'
+ ua = '-2.8887e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_9'
+ ub = '2.8956e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_9'
+ uc = 6.093e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0028+sky130_fd_pr__pfet_01v8_lvt__u0_diff_9'
+ a0 = '1.7177+sky130_fd_pr__pfet_01v8_lvt__a0_diff_9'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_9'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.20801+sky130_fd_pr__pfet_01v8_lvt__ags_diff_9'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_9'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_9'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_9+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0032329
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.027556
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9'
+ kt2 = -0.055045
+ at = 272010.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.425+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_10'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10'
+ ua = '-2.8587e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_10'
+ ub = '2.8956e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_10'
+ uc = 6.093e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0029+sky130_fd_pr__pfet_01v8_lvt__u0_diff_10'
+ a0 = '1.6516+sky130_fd_pr__pfet_01v8_lvt__a0_diff_10'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_10'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.2386+sky130_fd_pr__pfet_01v8_lvt__ags_diff_10'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_10'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_10'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_10+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0022476
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.020667
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.60135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10'
+ kt2 = -0.055045
+ at = 282740.0
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.35+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.04254+sky130_fd_pr__pfet_01v8_lvt__k2_diff_11'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '103960+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11'
+ ua = '-2.952e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_11'
+ ub = '3.2562e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_11'
+ uc = 5.0516e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0033729+sky130_fd_pr__pfet_01v8_lvt__u0_diff_11'
+ a0 = '1.494+sky130_fd_pr__pfet_01v8_lvt__a0_diff_11'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_11'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.3059+sky130_fd_pr__pfet_01v8_lvt__ags_diff_11'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_11'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_11'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_11+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '3.9645+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.097732
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.087651
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.65196+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11'
+ kt2 = -0.056015
+ at = 25215.0
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.39+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_12'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12'
+ ua = '-2.812e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_12'
+ ub = '2.9317e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_12'
+ uc = 6.4764e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0033729+sky130_fd_pr__pfet_01v8_lvt__u0_diff_12'
+ a0 = '1.494+sky130_fd_pr__pfet_01v8_lvt__a0_diff_12'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_12'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.3059+sky130_fd_pr__pfet_01v8_lvt__ags_diff_12'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_12'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_12'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_12+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '3.9645+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.043596
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.066402
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.65828+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12'
+ kt2 = -0.050974
+ at = 62896.0
+ ute = -0.43434
+ ua1 = 8.9635e-10
+ ub1 = -6.3517e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1.495e-06 lmax = 1.505e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.41071+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_13'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '70582+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13'
+ ua = '-3.0457e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_13'
+ ub = '3.1477e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_13'
+ uc = 6.9044e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0027+sky130_fd_pr__pfet_01v8_lvt__u0_diff_13'
+ a0 = '1.6213+sky130_fd_pr__pfet_01v8_lvt__a0_diff_13'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_13'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.55538+sky130_fd_pr__pfet_01v8_lvt__ags_diff_13'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_13'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_13'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_13+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.00979
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.032147
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13'
+ kt2 = -0.075412
+ at = 120290.0
+ ute = -0.13298
+ ua1 = 6.6751e-10
+ ub1 = -1.094e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.40571+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_14'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '128330+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14'
+ ua = '-3.0057e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_14'
+ ub = '3.1477e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_14'
+ uc = 7.5872e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0028528+sky130_fd_pr__pfet_01v8_lvt__u0_diff_14'
+ a0 = '1.4098+sky130_fd_pr__pfet_01v8_lvt__a0_diff_14'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_14'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.53402+sky130_fd_pr__pfet_01v8_lvt__ags_diff_14'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_14'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_14'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_14+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0178
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.042209
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.60135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14'
+ kt2 = -0.035779
+ at = 225860.0
+ ute = -0.17021
+ ua1 = 6.4145e-10
+ ub1 = -1.094e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 3.370e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.4+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_15'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15'
+ ua = '-3.0179e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_15'
+ ub = '3.0842e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_15'
+ uc = 5.6056e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0026+sky130_fd_pr__pfet_01v8_lvt__u0_diff_15'
+ a0 = '1.6516+sky130_fd_pr__pfet_01v8_lvt__a0_diff_15'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_15'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.4+sky130_fd_pr__pfet_01v8_lvt__ags_diff_15'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_15'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_15'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_15+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0068633
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.030692
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15'
+ kt2 = -0.055045
+ at = 247530.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.41+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_16'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16'
+ ua = '-2.9587e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_16'
+ ub = '2.9656e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_16'
+ uc = 4.8744e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0026+sky130_fd_pr__pfet_01v8_lvt__u0_diff_16'
+ a0 = '1.6516+sky130_fd_pr__pfet_01v8_lvt__a0_diff_16'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_16'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.32454+sky130_fd_pr__pfet_01v8_lvt__ags_diff_16'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_16'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_16'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_16+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0031348
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.022409
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16'
+ kt2 = -0.055045
+ at = 272010.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.425+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_17'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17'
+ ua = '-2.9587e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_17'
+ ub = '2.9656e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_17'
+ uc = 4.8744e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0026+sky130_fd_pr__pfet_01v8_lvt__u0_diff_17'
+ a0 = '1.6516+sky130_fd_pr__pfet_01v8_lvt__a0_diff_17'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_17'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.26919+sky130_fd_pr__pfet_01v8_lvt__ags_diff_17'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_17'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_17'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_17+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0016443
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.0177
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.60135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17'
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.37557+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_18'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '96388+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18'
+ ua = '-2.8839e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_18'
+ ub = '3.162e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_18'
+ uc = 6.3138e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0035466+sky130_fd_pr__pfet_01v8_lvt__u0_diff_18'
+ a0 = '1+sky130_fd_pr__pfet_01v8_lvt__a0_diff_18'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_18'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.42941+sky130_fd_pr__pfet_01v8_lvt__ags_diff_18'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_18'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_18'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_18+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.099935
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.065849
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62196+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18'
+ kt2 = -0.056015
+ at = 25215.0
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.385+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_19'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '182010+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19'
+ ua = '-2.8124e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_19'
+ ub = '2.9317e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_19'
+ uc = 6.0062e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0033+sky130_fd_pr__pfet_01v8_lvt__u0_diff_19'
+ a0 = '1.6516+sky130_fd_pr__pfet_01v8_lvt__a0_diff_19'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_19'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.3408+sky130_fd_pr__pfet_01v8_lvt__ags_diff_19'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_19'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_19'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_19+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.051183
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.056281
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.63828+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19'
+ kt2 = -0.056015
+ at = 59336.0
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1.495e-06 lmax = 1.505e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.41857+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_20'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '90748+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20'
+ ua = '-2.9616e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_20'
+ ub = '3.029e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_20'
+ uc = 7.1536e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00285+sky130_fd_pr__pfet_01v8_lvt__u0_diff_20'
+ a0 = '1+sky130_fd_pr__pfet_01v8_lvt__a0_diff_20'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_20'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.26966+sky130_fd_pr__pfet_01v8_lvt__ags_diff_20'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_20'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_20'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_20+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.010422
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.025214
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20'
+ kt2 = -0.055045
+ at = 152260.0
+ ute = -0.13298
+ ua1 = 6.6129e-10
+ ub1 = -1.094e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.42357+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.054915+sky130_fd_pr__pfet_01v8_lvt__k2_diff_21'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '91111+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21'
+ ua = '-2.8653e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_21'
+ ub = '2.9727e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_21'
+ uc = '7.2624e-011+sky130_fd_pr__pfet_01v8_lvt__uc_diff_21'
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00325+sky130_fd_pr__pfet_01v8_lvt__u0_diff_21'
+ a0 = '1.064+sky130_fd_pr__pfet_01v8_lvt__a0_diff_21'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_21'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.47558+sky130_fd_pr__pfet_01v8_lvt__ags_diff_21'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_21'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_21'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.19645+sky130_fd_pr__pfet_01v8_lvt__voff_diff_21+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5069+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.015362
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.032745
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.56135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21'
+ kt2 = -0.035779
+ at = 126070.0
+ ute = -0.22808
+ ua1 = 6.6129e-10
+ ub1 = -1.1159e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.41857+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_22'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '90748+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22'
+ ua = '-2.7794e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_22'
+ ub = '2.7289e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_22'
+ uc = '6.0493e-011+sky130_fd_pr__pfet_01v8_lvt__uc_diff_22'
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0029012+sky130_fd_pr__pfet_01v8_lvt__u0_diff_22'
+ a0 = '1+sky130_fd_pr__pfet_01v8_lvt__a0_diff_22'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_22'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.16045+sky130_fd_pr__pfet_01v8_lvt__ags_diff_22'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_22'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_22'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_22+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0069872
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.023147
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22'
+ kt2 = -0.055045
+ at = 165690.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -8.6535e-20
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.42+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_23'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23'
+ ua = '-2.9465e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_23'
+ ub = '2.9527e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_23'
+ uc = 6.093e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0026321+sky130_fd_pr__pfet_01v8_lvt__u0_diff_23'
+ a0 = '1.5459+sky130_fd_pr__pfet_01v8_lvt__a0_diff_23'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_23'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.35163+sky130_fd_pr__pfet_01v8_lvt__ags_diff_23'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_23'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_23'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_23+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0036208
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.021411
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.59135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23'
+ kt2 = -0.055045
+ at = 272010.0
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.42+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_24'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24'
+ ua = '-3.0054e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_24'
+ ub = '3.0419e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_24'
+ uc = 4.9353e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.002524+sky130_fd_pr__pfet_01v8_lvt__u0_diff_24'
+ a0 = '1.6387+sky130_fd_pr__pfet_01v8_lvt__a0_diff_24'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_24'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.31668+sky130_fd_pr__pfet_01v8_lvt__ags_diff_24'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_24'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_24'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_24+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.60135+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24'
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.37557+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_25'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '91569+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25'
+ ua = '-2.8839e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_25'
+ ub = '3.162e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_25'
+ uc = 6.3138e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0035466+sky130_fd_pr__pfet_01v8_lvt__u0_diff_25'
+ a0 = '1+sky130_fd_pr__pfet_01v8_lvt__a0_diff_25'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_25'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.42512+sky130_fd_pr__pfet_01v8_lvt__ags_diff_25'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_25'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_25'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_25+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.11592
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.052679
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.62196+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25'
+ kt2 = -0.056015
+ at = 25215.0
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.41757+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.048341+sky130_fd_pr__pfet_01v8_lvt__k2_diff_26'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '107140+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26'
+ ua = '-2.9416e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_26'
+ ub = '3.122e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_26'
+ uc = 6.9452e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00325+sky130_fd_pr__pfet_01v8_lvt__u0_diff_26'
+ a0 = '1+sky130_fd_pr__pfet_01v8_lvt__a0_diff_26'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_26'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.42087+sky130_fd_pr__pfet_01v8_lvt__ags_diff_26'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_26'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_26'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_26+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.053903
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.04425
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.63196+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26'
+ kt2 = -0.056015
+ at = 59336.0
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.29+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.032091+sky130_fd_pr__pfet_01v8_lvt__k2_diff_27'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27'
+ ua = '-2.7692e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_27'
+ ub = '2.877e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_27'
+ uc = 7.4772e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00284+sky130_fd_pr__pfet_01v8_lvt__u0_diff_27'
+ a0 = '1.2885+sky130_fd_pr__pfet_01v8_lvt__a0_diff_27'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_27'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_27'
+ b0 = '-2.8192e-008+sky130_fd_pr__pfet_01v8_lvt__b0_diff_27'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_27'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_27+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.18497+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.016674
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.030802
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.57503+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27'
+ kt2 = -0.085339
+ at = 191800.0
+ ute = -0.138
+ ua1 = 6.7978e-10
+ ub1 = -1.3904e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.385+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.024785+sky130_fd_pr__pfet_01v8_lvt__k2_diff_28'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28'
+ ua = '-2.9266e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_28'
+ ub = '2.8835e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_28'
+ uc = 6.0125e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0024126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_28'
+ a0 = '1.6218+sky130_fd_pr__pfet_01v8_lvt__a0_diff_28'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_28'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_28'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_28'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_28'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_28+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.18497+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.00013293
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01462
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.61455+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28'
+ kt2 = -0.055045
+ at = 290160.0
+ ute = -0.17727
+ ua1 = 6.8217e-10
+ ub1 = -1.7565e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.365+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.024785+sky130_fd_pr__pfet_01v8_lvt__k2_diff_29'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29'
+ ua = '-2.9966e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_29'
+ ub = '3.035e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_29'
+ uc = 6.6138e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0025126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_29'
+ a0 = '1.4529+sky130_fd_pr__pfet_01v8_lvt__a0_diff_29'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_29'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.20729+sky130_fd_pr__pfet_01v8_lvt__ags_diff_29'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_29'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_29'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_29+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.18497+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0076315
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.023279
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.600+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29'
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -0.11107
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.35+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.024785+sky130_fd_pr__pfet_01v8_lvt__k2_diff_30'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30'
+ ua = '-2.9966e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_30'
+ ub = '3.035e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_30'
+ uc = 6.6138e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0024126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_30'
+ a0 = '1.5205+sky130_fd_pr__pfet_01v8_lvt__a0_diff_30'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_30'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_30'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_30'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_30'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_30+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.18497+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0058704
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.027069
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.61457+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30'
+ kt2 = -0.055045
+ at = 269260.0
+ ute = -0.095746
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.375+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.024785+sky130_fd_pr__pfet_01v8_lvt__k2_diff_31'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31'
+ ua = '-2.9266e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_31'
+ ub = '2.8835e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_31'
+ uc = 6.0125e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0024126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_31'
+ a0 = '1.4529+sky130_fd_pr__pfet_01v8_lvt__a0_diff_31'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_31'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_31'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_31'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_31'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_31+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.18497+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.001223
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.020201
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.61455+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31'
+ kt2 = -0.055045
+ at = 273740.0
+ ute = -0.17727
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.35+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.015793+sky130_fd_pr__pfet_01v8_lvt__k2_diff_32'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '101480+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32'
+ ua = '-3.01e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_32'
+ ub = '3.2578e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_32'
+ uc = 6.5372e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0028126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_32'
+ a0 = '1.6894+sky130_fd_pr__pfet_01v8_lvt__a0_diff_32'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_32'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_32'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_32'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_32'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_32+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.06289+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.098214
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.079955
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.63756+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32'
+ kt2 = -0.085339
+ at = 10582.0
+ ute = -0.21235
+ ua1 = 7.2317e-10
+ ub1 = -2.3247e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.307+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.015793+sky130_fd_pr__pfet_01v8_lvt__k2_diff_33'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '168310+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33'
+ ua = '-2.9492e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_33'
+ ub = '3.1278e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_33'
+ uc = 7.4286e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0029126+sky130_fd_pr__pfet_01v8_lvt__u0_diff_33'
+ a0 = '1.6894+sky130_fd_pr__pfet_01v8_lvt__a0_diff_33'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_33'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.15242+sky130_fd_pr__pfet_01v8_lvt__ags_diff_33'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_33'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_33'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_33+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.06289+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.041068
+ pdiblcb = -0.025
+ drout = 0.42626
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.054764
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.57831+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33'
+ kt2 = -0.085339
+ at = 126490.0
+ ute = -0.1
+ ua1 = 6.9424e-10
+ ub1 = -1.0948e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.3585+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.036577+sky130_fd_pr__pfet_01v8_lvt__k2_diff_34'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '93472+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34'
+ ua = '-2.7682e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_34'
+ ub = '2.7913e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_34'
+ uc = 7.3044e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.002898+sky130_fd_pr__pfet_01v8_lvt__u0_diff_34'
+ a0 = '1.3185+sky130_fd_pr__pfet_01v8_lvt__a0_diff_34'
+ keta = '-0.011825+sky130_fd_pr__pfet_01v8_lvt__keta_diff_34'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.47+sky130_fd_pr__pfet_01v8_lvt__ags_diff_34'
+ b0 = '4.9905e-008+sky130_fd_pr__pfet_01v8_lvt__b0_diff_34'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_34'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_34+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.020189
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.031365
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.57819+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34'
+ kt2 = -0.085339
+ at = 110630.0
+ ute = -0.1
+ ua1 = 7.2317e-10
+ ub1 = -9.3948e-20
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.33+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.037416+sky130_fd_pr__pfet_01v8_lvt__k2_diff_35'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35'
+ ua = '-3.0809e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_35'
+ ub = '3.1278e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_35'
+ uc = 5.4659e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00217+sky130_fd_pr__pfet_01v8_lvt__u0_diff_35'
+ a0 = '1.6894+sky130_fd_pr__pfet_01v8_lvt__a0_diff_35'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_35'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.31912+sky130_fd_pr__pfet_01v8_lvt__ags_diff_35'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_35'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_35'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_35+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0071618
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.024552
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.64457+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35'
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -0.095746
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.34+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.037416+sky130_fd_pr__pfet_01v8_lvt__k2_diff_36'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36'
+ ua = '-3.0709e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_36'
+ ub = '3.1078e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_36'
+ uc = 5.4659e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.002166+sky130_fd_pr__pfet_01v8_lvt__u0_diff_36'
+ a0 = '1.6894+sky130_fd_pr__pfet_01v8_lvt__a0_diff_36'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_36'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.23815+sky130_fd_pr__pfet_01v8_lvt__ags_diff_36'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_36'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_36'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_36+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0030771
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.018053
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.64457+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36'
+ kt2 = -0.055045
+ at = 269260.0
+ ute = -0.095746
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.36+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.037416+sky130_fd_pr__pfet_01v8_lvt__k2_diff_37'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '123760+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37'
+ ua = '-3.0306e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_37'
+ ub = '3.077e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_37'
+ uc = 6.0065e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.00228+sky130_fd_pr__pfet_01v8_lvt__u0_diff_37'
+ a0 = '1.7239+sky130_fd_pr__pfet_01v8_lvt__a0_diff_37'
+ keta = '-0.01258+sky130_fd_pr__pfet_01v8_lvt__keta_diff_37'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.26461+sky130_fd_pr__pfet_01v8_lvt__ags_diff_37'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_37'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_37'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_37+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.00043292
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.013574
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.67455+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37'
+ kt2 = -0.055045
+ at = 282210.0
+ ute = -0.28592
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos
* DC IV MOS Parameters
+ lmin = 3.45e-07 lmax = 3.55e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.2655+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.016213+sky130_fd_pr__pfet_01v8_lvt__k2_diff_38'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '74652+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38'
+ ua = '-3.0256e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_38'
+ ub = '3.3481e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_38'
+ uc = 5.7404e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0027427+sky130_fd_pr__pfet_01v8_lvt__u0_diff_38'
+ a0 = '1.1627+sky130_fd_pr__pfet_01v8_lvt__a0_diff_38'
+ keta = '-0.011825+sky130_fd_pr__pfet_01v8_lvt__keta_diff_38'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.23897+sky130_fd_pr__pfet_01v8_lvt__ags_diff_38'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_38'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_38'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_38+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.14839
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.037022
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.63756+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38'
+ kt2 = -0.085339
+ at = 10582.0
+ ute = -0.21235
+ ua1 = 7.2317e-10
+ ub1 = -2.3247e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = '2.8e-009+sky130_fd_pr__pfet_01v8_lvt__lint_diff'
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = '7.476e-009+sky130_fd_pr__pfet_01v8_lvt__wint_diff'
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = '4.23e-009*sky130_fd_pr__pfet_01v8_lvt__toxe_mult+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8_lvt__toxe_mult*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))'
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = '1*sky130_fd_pr__pfet_01v8_lvt__rshp_mult'
* Threshold Voltage Parameters
+ vth0 = '-0.2655+sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))'
+ k1 = 0.64774
+ k2 = '-0.016213+sky130_fd_pr__pfet_01v8_lvt__k2_diff_39'
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = '96343+sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39'
+ ua = '-2.9058e-009+sky130_fd_pr__pfet_01v8_lvt__ua_diff_39'
+ ub = '3.0795e-018+sky130_fd_pr__pfet_01v8_lvt__ub_diff_39'
+ uc = 6.7633e-11
+ rdsw = '484.7+sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39'
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = '0.0025803+sky130_fd_pr__pfet_01v8_lvt__u0_diff_39'
+ a0 = '1.1627+sky130_fd_pr__pfet_01v8_lvt__a0_diff_39'
+ keta = '-0.011825+sky130_fd_pr__pfet_01v8_lvt__keta_diff_39'
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = '0.5+sky130_fd_pr__pfet_01v8_lvt__ags_diff_39'
+ b0 = '0+sky130_fd_pr__pfet_01v8_lvt__b0_diff_39'
+ b1 = '2.1073e-024+sky130_fd_pr__pfet_01v8_lvt__b1_diff_39'
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = '-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_diff_39+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))'
+ nfactor = '2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))'
+ tvoff = '0+sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39'
+ tvfbsdoff = 0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 0.0001
+ cdscd = 1.0e-10
+ eta0 = '0.2+sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39'
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = '0.030097+sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39'
+ pdiblc1 = 0.0
+ pdiblc2 = 0.077088
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.034486
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = '0+sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39'
+ pditsl = 0.0
+ pditsd = '0+sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39'
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = '0+sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39'
+ bgidl = '2.3e009+sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39'
+ cgidl = '0.5+sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39'
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = '-0.61219+sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39'
+ kt2 = -0.085339
+ at = 100240.0
+ ute = -0.10000
+ ua1 = 7.2317e-10
+ ub1 = -2.7896e-19
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgso = '1e-010*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cgdl = '0*sky130_fd_pr__pfet_01v8_lvt__overlap_mult'
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = '0+sky130_fd_pr__pfet_01v8_lvt__dlc_diff+sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak'
+ dwc = '0+sky130_fd_pr__pfet_01v8_lvt__dwc_diff'
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = '0.00076823*sky130_fd_pr__pfet_01v8_lvt__ajunction_mult'
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = '9.152e-011*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = '2.3894e-010*sky130_fd_pr__pfet_01v8_lvt__pjunction_mult'
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = '0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff'
+ kvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff'
+ lkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff'
+ wkvth0 = '0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff'
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = '0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff'
+ lku0 = '0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff'
+ wku0 = '0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff'
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = '0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff'
+ steta0 = 0.0
+ tku0 = 0.0
.ends pfet_01v8_lvt
