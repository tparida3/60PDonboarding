* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.model diode_pw2nd_05v5 d
+ level = 3.0
+ tlevc = 1.0
+ area = 1.0e+12
* Junction Capacitance Parameters
+ cj = '0.0013459*1e-12*sky130_fd_pr__nfet_01v8__ajunction_mult' $ Units: farad/meter^2
+ mj = 0.44
+ pb = 0.729 $ Units: volt
+ cjsw = '3.6001e-011*1e-6*sky130_fd_pr__nfet_01v8__pjunction_mult' $ Units: farad/meter
+ mjsw = 0.0009
+ php = 0.2 $ Units: volt
+ cta = 0.000792 $ Units: 1/coulomb
+ ctp = 1e-005 $ Units: 1/coulomb
+ tpb = 0.0012287 $ Units: volt/coulomb
+ tphp = 0 $ Units: volt/coulomb
* Diode IV Parameters
+ js = 2.75e-015 $ Units: amper/meter^2
+ jsw = 6e-016 $ Units: amper/meter
+ n = 1.2928
+ rs = 981 $ Units: ohm (ohm/meter^2 if area defined)
+ ik = '1.3e-009/1e-12' $ Units: amper/meter^2
+ ikr = '0/1e-12' $ Units: amper/meter^2
+ vb = 11.7 $ Units: volt
+ ibv = 0.00106 $ Units: amper
+ trs = 0 $ Units: 1/coulomb
+ eg = 1.05 $ Units: electron-volt
+ xti = 2.0
+ tref = 30 $ Units: coulomb
* Default Parameters
+ tcv = 0 $ Units: 1/coulomb
+ gap1 = 0.000473 $ Units: electron-volt/coulomb
+ gap2 = 1110.0
+ ttt1 = 0 $ Units: 1/coulomb
+ ttt2 = 0 $ Units: 1/coulomb^2
+ tm1 = 0 $ Units: 1/coulomb
+ tm2 = 0 $ Units: 1/coulomb^2
+ lm = 0 $ Units: meter
+ lp = 0 $ Units: meter
+ wm = 0 $ Units: meter
+ wp = 0 $ Units: meter
+ xm = 0 $ Units: meter
+ xoi = 10000.0
+ xom = 10000 $ Units: angstrom
+ xp = 0 $ Units: meter
+ xw = 0 $ Units: meter
